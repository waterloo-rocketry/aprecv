module srad_aprs_receiver_tb;
endmodule
