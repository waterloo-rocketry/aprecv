module filter_iir #(
) (
);

endmodule
