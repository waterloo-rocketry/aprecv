module srad_aprs_receiver_top;
endmodule
